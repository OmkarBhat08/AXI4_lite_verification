`define ADDR_WIDTH 4
`define DATA_WIDTH 32
