class base_seq extends uvm_sequence #(axi4_seq_item);
  `uvm_object_utils(base_seq)
  
  function new(string name="base_seq"); 
    super.new(name); 
  endfunction
  
  task body();
    axi4_seq_item req;
    `uvm_info(get_type_name(), " ------ Base Sequence ------ ", UVM_LOW)
    repeat (3) begin
      req = axi4_seq_item::type_id::create("req");
      start_item(req);
      assert(req.randomize() with { req.BREADY == 1;} );
      finish_item(req);
    end
  endtask
endclass

// -----------------------------------------------------------------
// Simple write with strobe = 'b1111
class simple_write extends base_seq;
  `uvm_object_utils(simple_write)

  function new(string name = "simple_write");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Simple write with strobe = 'b1111 ------ ", UVM_LOW)
    repeat(1) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.AWADDR inside {0}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.AWADDR inside {4}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.AWADDR inside {8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Simple read
class simple_read extends base_seq;
  `uvm_object_utils(simple_read)

  function new(string name = "simple_read");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Simple read ------ ", UVM_LOW)
    repeat(3) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.ARADDR inside {0, 4, 8}; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})

    end
  endtask
endclass

// -----------------------------------------------------------------
// Read followed by Write
class read_followed_by_write extends base_seq;
  `uvm_object_utils(read_followed_by_write)
  bit [`ADDR_WIDTH-1:0] prev_addr;

  function new(string name = "read_followed_by_write");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Read followed by Write ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WSTRB == 4'b1111; req.WVALID == 1; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.AWADDR == prev_addr; req.AWVALID == 0; req.WSTRB == 4'b1111; req.WVALID == 0; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Parallel Read and Write
class parallel_read_write extends base_seq;
  `uvm_object_utils(parallel_read_write)

  function new(string name = "parallel_read_write");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Parallel Read and Write ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WSTRB == 4'b1111; req.WVALID == 1; req.ARADDR inside {0,4,8}; req.ARVALID == 1; req.RREADY == 1;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Write data before address
class data_before_addr extends base_seq;
  `uvm_object_utils(data_before_addr)

  function new(string name = "data_before_addr");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Write data before address ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.ARVALID == 0; req.RREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Write address before data together
class addr_before_data extends base_seq;
  `uvm_object_utils(addr_before_data)

  function new(string name = "addr_before_data");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Write address before data together ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.ARVALID == 0; req.RREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Write address and data together
class data_with_addr extends base_seq;
  `uvm_object_utils(data_with_addr)

  function new(string name = "data_with_addr");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Write address and data together ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.ARVALID == 0; req.RREADY == 0; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Back to back write to same address and read
class continuous_write extends base_seq;
  `uvm_object_utils(continuous_write)
  bit [`ADDR_WIDTH-1:0] prev_addr;
  bit [`DATA_WIDTH-1:0] prev_data;

  function new(string name = "continuous_write");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Back to back write to same address and read ------ ", UVM_LOW)
    prev_addr = 0;
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR != prev_addr; req.AWVALID == 1; req.WSTRB == 4'b1111; req.WVALID == 1; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      prev_data = req.WDATA;

      `uvm_do_with(req, {req.AWADDR == prev_addr; req.AWVALID == 1; req.WSTRB == 4'b1111; req.WVALID == 1; req.WDATA != prev_data; req.ARVALID == 0; req.RREADY == 0;})
      prev_data = req.WDATA;

      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Write with strobe select and read back from the same address
class write_strobe_select_1 extends base_seq;
  `uvm_object_utils(write_strobe_select_1)
  bit [`ADDR_WIDTH-1:0] prev_addr;

  function new(string name = "write_strobe_select_1");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Write with strobe select and read back from the same address  ------ ", UVM_LOW)
    repeat(3) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB inside {[0:15]}; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
    end
  endtask
endclass

class write_strobe_select_2 extends base_seq;
  `uvm_object_utils(write_strobe_select_2)
  bit [`ADDR_WIDTH-1:0] prev_addr;

  function new(string name = "write_strobe_select_2");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Write with strobe select and read back from the same address  ------ ", UVM_LOW)
    repeat(3) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b0001; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})

      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b0010; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})

      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b0100; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})

      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1000; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// BVALID Hold
class bvalid_hold_seq extends base_seq;
  `uvm_object_utils(bvalid_hold_seq)
  bit [`ADDR_WIDTH-1:0] prev_addr;

  function new(string name = "bvalid_hold_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), $sformatf(" ------ BVALID Hold ------ "), UVM_LOW)
    repeat(5) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.BREADY == 0; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.AWADDR == prev_addr; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.BREADY == 0; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.AWADDR == prev_addr; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.BREADY == 0; req.ARVALID == 0; req.RREADY == 0;})
      `uvm_do_with(req, {req.AWADDR == prev_addr; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.ARVALID == 0; req.RREADY == 0;})
    end
  endtask
endclass
// -----------------------------------------------------------------
// RVALID Hold
class rvalid_hold_seq extends base_seq;
  `uvm_object_utils(rvalid_hold_seq)
  bit [`ADDR_WIDTH-1:0] prev_addr;

  function new(string name = "rvalid_hold_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), $sformatf(" ------ BVALID Hold ------ "), UVM_LOW)
    repeat(5) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111; req.BREADY == 0; req.ARVALID == 0; req.RREADY == 0;})
      prev_addr = req.AWADDR;
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 0; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 0; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 0; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
      `uvm_do_with(req, {req.ARADDR == prev_addr; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Invalid Address Write and Read

class invalid_addr extends base_seq;
  `uvm_object_utils(invalid_addr)

  function new(string name = "invalid_addr");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), $sformatf(" ------ invalid address write and read ------ "), UVM_LOW)
    repeat(10) begin
      req = axi4_seq_item::type_id::create("req");
      `uvm_do_with(req, {req.ARVALID == 1; req.RREADY == 1; req.AWADDR inside {0,4,8}; req.AWVALID == 1; req.WVALID == 1; req.WSTRB == 4'b1111;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Interrupt High
class irq_seq_1 extends base_seq;
  `uvm_object_utils(irq_seq_1)

  function new(string name = "irq_seq_1");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), $sformatf(" ------ Interrupt High ------ "), UVM_LOW)
    repeat(2) begin
      `uvm_do_with(req, {req.AWADDR == 8; req.AWVALID == 1; req.WSTRB[0] == 1; req.WDATA[0] == 1; req.WVALID == 1; req.EXT_IRQ_IN == 1;})
      #1000000;
      `uvm_do_with(req, {req.ARADDR == 8; req.ARVALID == 1; req.RREADY == 1; req.AWVALID == 0; req.WVALID == 0; req.BREADY == 0; req.EXT_IRQ_IN == 1;})
    end
  endtask
endclass

// -----------------------------------------------------------------
// Interrupt 

class irq_seq_2 extends base_seq;
  `uvm_object_utils(irq_seq_2)

  function new(string name = "irq_seq_2");
    super.new(name);
  endfunction

  task body();
    `uvm_info(get_type_name(), " ------ Interrupt High ------ ", UVM_LOW)
    repeat(3) begin
      `uvm_do_with(req, {req.AWADDR == 8; req.AWVALID == 1; req.WSTRB[0] == 1; req.WDATA[0] == 1; req.WVALID == 1; req.EXT_IRQ_IN == 1;})
      #10_000;
      `uvm_do_with(req, {req.AWADDR == 8; req.AWVALID == 1; req.WSTRB[0] == 1; req.WDATA[0] == 1; req.WVALID == 1; req.EXT_IRQ_IN == 0;})
    end
  endtask
endclass

// -----------------------------------------------------------------

